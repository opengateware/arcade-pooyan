-- -----------------------------------------------------------------------
--
-- Syntiac's generic VHDL support files.
--
-- -----------------------------------------------------------------------
-- Copyright 2005-2008 by Peter Wendrich (pwsoft@syntiac.com)
-- http://www.syntiac.com/fpga64.html
--
-- Modified April 2016 by Dar (darfpga@aol.fr) 
-- http://darfpga.blogspot.fr
--   Remove address register when writing
--
-- -----------------------------------------------------------------------
--
-- gen_rwram.vhd
--
-- -----------------------------------------------------------------------
--
-- generic ram.
--
-- -----------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;

-- -----------------------------------------------------------------------

entity gen_ram is
    generic (
        dWidth : integer := 8;
        aWidth : integer := 10
    );
    port (
        clk  : in std_logic;
        we   : in std_logic;
        addr : in std_logic_vector((aWidth - 1) downto 0);
        d    : in std_logic_vector((dWidth - 1) downto 0);
        q    : out std_logic_vector((dWidth - 1) downto 0)
    );
end entity;

-- -----------------------------------------------------------------------

architecture rtl of gen_ram is
    subtype addressRange is integer range 0 to ((2 ** aWidth) - 1);
    type ramDef is array(addressRange) of std_logic_vector((dWidth - 1) downto 0);
    signal ram : ramDef;

    signal rAddrReg : std_logic_vector((aWidth - 1) downto 0);
    signal qReg : std_logic_vector((dWidth - 1) downto 0);
begin

    -- -----------------------------------------------------------------------
    -- Memory write
    -- -----------------------------------------------------------------------
    process (clk)
    begin
        if rising_edge(clk) then
            if we = '1' then
                ram(to_integer(unsigned(addr))) <= d;
            end if;
        end if;
    end process;

    -- -----------------------------------------------------------------------
    -- Memory read
    -- -----------------------------------------------------------------------
    process (clk)
    begin
        if rising_edge(clk) then
            q <= ram(to_integer(unsigned(addr)));
        end if;
    end process;

end architecture;
